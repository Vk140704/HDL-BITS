Implement the following circuit:
in----------out
  Answer 
module top_module (
    input in,
    output out);
wire w1;
    assign w1= in;
    assign out = w1;
endmodule

